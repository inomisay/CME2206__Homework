library verilog;
use verilog.vl_types.all;
entity Yasamin_2022510013_Group31_ALU_vlg_check_tst is
    port(
        OUTPUT          : in     vl_logic_vector(3 downto 0);
        Overflow        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Yasamin_2022510013_Group31_ALU_vlg_check_tst;
